module our_OnOff(
	input a,
	input b,
	output c
);

	assign c = a ^ b;
endmodule
